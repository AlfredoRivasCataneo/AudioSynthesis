library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity EnvelopeGenerator is
end EnvelopeGenerator;

architecture Behavioral of EnvelopeGenerator is

begin


end Behavioral;

