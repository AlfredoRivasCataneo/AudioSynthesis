library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
entity sinewave is
port (clksen :in  std_logic;
dataout : out std_logic_vector(15 downto 0);
);
end sinewave;
architecture Behavioral of SineWave is


constant D0: std_logic_vector(15 downto 0) := x"80";
constant D1: std_logic_vector(15 downto 0) := x"82";
constant D2: std_logic_vector(15 downto 0) := x"84";
constant D3: std_logic_vector(15 downto 0) := x"87";
constant D4: std_logic_vector(15 downto 0) := x"89";
constant D5: std_logic_vector(15 downto 0) := x"8B";
constant D6: std_logic_vector(15 downto 0) := x"8D";
constant D7: std_logic_vector(15 downto 0) := x"90";
constant D8: std_logic_vector(15 downto 0) := x"92";
constant D9: std_logic_vector(15 downto 0) := x"94";
constant D10: std_logic_vector(15 downto 0) := x"96";
constant D11: std_logic_vector(15 downto 0) := x"98";
constant D12: std_logic_vector(15 downto 0) := x"9B";
constant D13: std_logic_vector(15 downto 0) := x"9D";
constant D14: std_logic_vector(15 downto 0) := x"9F";
constant D15: std_logic_vector(15 downto 0) := x"A1";
constant D16: std_logic_vector(15 downto 0) := x"A3";
constant D17: std_logic_vector(15 downto 0) := x"A5";
constant D18: std_logic_vector(15 downto 0) := x"A8";
constant D19: std_logic_vector(15 downto 0) := x"AA";
constant D20: std_logic_vector(15 downto 0) := x"AC";
constant D21: std_logic_vector(15 downto 0) := x"AE";
constant D22: std_logic_vector(15 downto 0) := x"B0";
constant D23: std_logic_vector(15 downto 0) := x"B2";
constant D24: std_logic_vector(15 downto 0) := x"B4";
constant D25: std_logic_vector(15 downto 0) := x"B6";
constant D26: std_logic_vector(15 downto 0) := x"B8";
constant D27: std_logic_vector(15 downto 0) := x"BA";
constant D28: std_logic_vector(15 downto 0) := x"BC";
constant D29: std_logic_vector(15 downto 0) := x"BE";
constant D30: std_logic_vector(15 downto 0) := x"C0";
constant D31: std_logic_vector(15 downto 0) := x"C2";
constant D32: std_logic_vector(15 downto 0) := x"C4";
constant D33: std_logic_vector(15 downto 0) := x"C6";
constant D34: std_logic_vector(15 downto 0) := x"C8";
constant D35: std_logic_vector(15 downto 0) := x"C9";
constant D36: std_logic_vector(15 downto 0) := x"CB";
constant D37: std_logic_vector(15 downto 0) := x"CD";
constant D38: std_logic_vector(15 downto 0) := x"CF";
constant D39: std_logic_vector(15 downto 0) := x"D1";
constant D40: std_logic_vector(15 downto 0) := x"D2";
constant D41: std_logic_vector(15 downto 0) := x"D4";
constant D42: std_logic_vector(15 downto 0) := x"D6";
constant D43: std_logic_vector(15 downto 0) := x"D7";
constant D44: std_logic_vector(15 downto 0) := x"D9";
constant D45: std_logic_vector(15 downto 0) := x"DB";
constant D46: std_logic_vector(15 downto 0) := x"DC";
constant D47: std_logic_vector(15 downto 0) := x"DE";
constant D48: std_logic_vector(15 downto 0) := x"DF";
constant D49: std_logic_vector(15 downto 0) := x"E1";
constant D50: std_logic_vector(15 downto 0) := x"E2";
constant D51: std_logic_vector(15 downto 0) := x"E3";
constant D52: std_logic_vector(15 downto 0) := x"E5";
constant D53: std_logic_vector(15 downto 0) := x"E6";
constant D54: std_logic_vector(15 downto 0) := x"E8";
constant D55: std_logic_vector(15 downto 0) := x"E9";
constant D56: std_logic_vector(15 downto 0) := x"EA";
constant D57: std_logic_vector(15 downto 0) := x"EB";
constant D58: std_logic_vector(15 downto 0) := x"ED";
constant D59: std_logic_vector(15 downto 0) := x"EE";
constant D60: std_logic_vector(15 downto 0) := x"EF";
constant D61: std_logic_vector(15 downto 0) := x"F0";
constant D62: std_logic_vector(15 downto 0) := x"F1";
constant D63: std_logic_vector(15 downto 0) := x"F2";
constant D64: std_logic_vector(15 downto 0) := x"F3";
constant D65: std_logic_vector(15 downto 0) := x"F4";
constant D66: std_logic_vector(15 downto 0) := x"F5";
constant D67: std_logic_vector(15 downto 0) := x"F6";
constant D68: std_logic_vector(15 downto 0) := x"F7";
constant D69: std_logic_vector(15 downto 0) := x"F7";
constant D70: std_logic_vector(15 downto 0) := x"F8";
constant D71: std_logic_vector(15 downto 0) := x"F9";
constant D72: std_logic_vector(15 downto 0) := x"FA";
constant D73: std_logic_vector(15 downto 0) := x"FA";
constant D74: std_logic_vector(15 downto 0) := x"FB";
constant D75: std_logic_vector(15 downto 0) := x"FC";
constant D76: std_logic_vector(15 downto 0) := x"FC";
constant D77: std_logic_vector(15 downto 0) := x"FD";
constant D78: std_logic_vector(15 downto 0) := x"FD";
constant D79: std_logic_vector(15 downto 0) := x"FE";
constant D80: std_logic_vector(15 downto 0) := x"FE";
constant D81: std_logic_vector(15 downto 0) := x"FE";
constant D82: std_logic_vector(15 downto 0) := x"FF";
constant D83: std_logic_vector(15 downto 0) := x"FF";
constant D84: std_logic_vector(15 downto 0) := x"FF";
constant D85: std_logic_vector(15 downto 0) := x"FF";
constant D86: std_logic_vector(15 downto 0) := x"FF";
constant D87: std_logic_vector(15 downto 0) := x"FF";
constant D88: std_logic_vector(15 downto 0) := x"FF";
constant D89: std_logic_vector(15 downto 0) := x"FF";
constant D90: std_logic_vector(15 downto 0) := x"FF";
constant D91: std_logic_vector(15 downto 0) := x"FF";
constant D92: std_logic_vector(15 downto 0) := x"FF";
constant D93: std_logic_vector(15 downto 0) := x"FF";
constant D94: std_logic_vector(15 downto 0) := x"FF";
constant D95: std_logic_vector(15 downto 0) := x"FF";
constant D96: std_logic_vector(15 downto 0) := x"FF";
constant D97: std_logic_vector(15 downto 0) := x"FF";
constant D98: std_logic_vector(15 downto 0) := x"FF";
constant D99: std_logic_vector(15 downto 0) := x"FE";
constant D100: std_logic_vector(15 downto 0) := x"FE";
constant D101: std_logic_vector(15 downto 0) := x"FE";
constant D102: std_logic_vector(15 downto 0) := x"FD";
constant D103: std_logic_vector(15 downto 0) := x"FD";
constant D104: std_logic_vector(15 downto 0) := x"FC";
constant D105: std_logic_vector(15 downto 0) := x"FC";
constant D106: std_logic_vector(15 downto 0) := x"FB";
constant D107: std_logic_vector(15 downto 0) := x"FA";
constant D108: std_logic_vector(15 downto 0) := x"FA";
constant D109: std_logic_vector(15 downto 0) := x"F9";
constant D110: std_logic_vector(15 downto 0) := x"F8";
constant D111: std_logic_vector(15 downto 0) := x"F7";
constant D112: std_logic_vector(15 downto 0) := x"F7";
constant D113: std_logic_vector(15 downto 0) := x"F6";
constant D114: std_logic_vector(15 downto 0) := x"F5";
constant D115: std_logic_vector(15 downto 0) := x"F4";
constant D116: std_logic_vector(15 downto 0) := x"F3";
constant D117: std_logic_vector(15 downto 0) := x"F2";
constant D118: std_logic_vector(15 downto 0) := x"F1";
constant D119: std_logic_vector(15 downto 0) := x"F0";
constant D120: std_logic_vector(15 downto 0) := x"EF";
constant D121: std_logic_vector(15 downto 0) := x"EE";
constant D122: std_logic_vector(15 downto 0) := x"ED";
constant D123: std_logic_vector(15 downto 0) := x"EB";
constant D124: std_logic_vector(15 downto 0) := x"EA";
constant D125: std_logic_vector(15 downto 0) := x"E9";
constant D126: std_logic_vector(15 downto 0) := x"E8";
constant D127: std_logic_vector(15 downto 0) := x"E6";
constant D128: std_logic_vector(15 downto 0) := x"E5";
constant D129: std_logic_vector(15 downto 0) := x"E3";
constant D130: std_logic_vector(15 downto 0) := x"E2";
constant D131: std_logic_vector(15 downto 0) := x"E1";
constant D132: std_logic_vector(15 downto 0) := x"DF";
constant D133: std_logic_vector(15 downto 0) := x"DE";
constant D134: std_logic_vector(15 downto 0) := x"DC";
constant D135: std_logic_vector(15 downto 0) := x"DB";
constant D136: std_logic_vector(15 downto 0) := x"D9";
constant D137: std_logic_vector(15 downto 0) := x"D7";
constant D138: std_logic_vector(15 downto 0) := x"D6";
constant D139: std_logic_vector(15 downto 0) := x"D4";
constant D140: std_logic_vector(15 downto 0) := x"D2";
constant D141: std_logic_vector(15 downto 0) := x"D1";
constant D142: std_logic_vector(15 downto 0) := x"CF";
constant D143: std_logic_vector(15 downto 0) := x"CD";
constant D144: std_logic_vector(15 downto 0) := x"CB";
constant D145: std_logic_vector(15 downto 0) := x"C9";
constant D146: std_logic_vector(15 downto 0) := x"C8";
constant D147: std_logic_vector(15 downto 0) := x"C6";
constant D148: std_logic_vector(15 downto 0) := x"C4";
constant D149: std_logic_vector(15 downto 0) := x"C2";
constant D150: std_logic_vector(15 downto 0) := x"C0";
constant D151: std_logic_vector(15 downto 0) := x"BE";
constant D152: std_logic_vector(15 downto 0) := x"BC";
constant D153: std_logic_vector(15 downto 0) := x"BA";
constant D154: std_logic_vector(15 downto 0) := x"B8";
constant D155: std_logic_vector(15 downto 0) := x"B6";
constant D156: std_logic_vector(15 downto 0) := x"B4";
constant D157: std_logic_vector(15 downto 0) := x"B2";
constant D158: std_logic_vector(15 downto 0) := x"B0";
constant D159: std_logic_vector(15 downto 0) := x"AE";
constant D160: std_logic_vector(15 downto 0) := x"AC";
constant D161: std_logic_vector(15 downto 0) := x"AA";
constant D162: std_logic_vector(15 downto 0) := x"A8";
constant D163: std_logic_vector(15 downto 0) := x"A5";
constant D164: std_logic_vector(15 downto 0) := x"A3";
constant D165: std_logic_vector(15 downto 0) := x"A1";
constant D166: std_logic_vector(15 downto 0) := x"9F";
constant D167: std_logic_vector(15 downto 0) := x"9D";
constant D168: std_logic_vector(15 downto 0) := x"9B";
constant D169: std_logic_vector(15 downto 0) := x"98";
constant D170: std_logic_vector(15 downto 0) := x"96";
constant D171: std_logic_vector(15 downto 0) := x"94";
constant D172: std_logic_vector(15 downto 0) := x"92";
constant D173: std_logic_vector(15 downto 0) := x"90";
constant D174: std_logic_vector(15 downto 0) := x"8D";
constant D175: std_logic_vector(15 downto 0) := x"8B";
constant D176: std_logic_vector(15 downto 0) := x"89";
constant D177: std_logic_vector(15 downto 0) := x"87";
constant D178: std_logic_vector(15 downto 0) := x"84";
constant D179: std_logic_vector(15 downto 0) := x"82";
constant D180: std_logic_vector(15 downto 0) := x"80";
constant D181: std_logic_vector(15 downto 0) := x"7E";
constant D182: std_logic_vector(15 downto 0) := x"7C";
constant D183: std_logic_vector(15 downto 0) := x"79";
constant D184: std_logic_vector(15 downto 0) := x"77";
constant D185: std_logic_vector(15 downto 0) := x"75";
constant D186: std_logic_vector(15 downto 0) := x"73";
constant D187: std_logic_vector(15 downto 0) := x"70";
constant D188: std_logic_vector(15 downto 0) := x"6E";
constant D189: std_logic_vector(15 downto 0) := x"6C";
constant D190: std_logic_vector(15 downto 0) := x"6A";
constant D191: std_logic_vector(15 downto 0) := x"68";
constant D192: std_logic_vector(15 downto 0) := x"65";
constant D193: std_logic_vector(15 downto 0) := x"63";
constant D194: std_logic_vector(15 downto 0) := x"61";
constant D195: std_logic_vector(15 downto 0) := x"5F";
constant D196: std_logic_vector(15 downto 0) := x"5D";
constant D197: std_logic_vector(15 downto 0) := x"5B";
constant D198: std_logic_vector(15 downto 0) := x"58";
constant D199: std_logic_vector(15 downto 0) := x"56";
constant D200: std_logic_vector(15 downto 0) := x"54";
constant D201: std_logic_vector(15 downto 0) := x"52";
constant D202: std_logic_vector(15 downto 0) := x"50";
constant D203: std_logic_vector(15 downto 0) := x"4E";
constant D204: std_logic_vector(15 downto 0) := x"4C";
constant D205: std_logic_vector(15 downto 0) := x"4A";
constant D206: std_logic_vector(15 downto 0) := x"48";
constant D207: std_logic_vector(15 downto 0) := x"46";
constant D208: std_logic_vector(15 downto 0) := x"44";
constant D209: std_logic_vector(15 downto 0) := x"42";
constant D210: std_logic_vector(15 downto 0) := x"40";
constant D211: std_logic_vector(15 downto 0) := x"3E";
constant D212: std_logic_vector(15 downto 0) := x"3C";
constant D213: std_logic_vector(15 downto 0) := x"3A";
constant D214: std_logic_vector(15 downto 0) := x"38";
constant D215: std_logic_vector(15 downto 0) := x"37";
constant D216: std_logic_vector(15 downto 0) := x"35";
constant D217: std_logic_vector(15 downto 0) := x"33";
constant D218: std_logic_vector(15 downto 0) := x"31";
constant D219: std_logic_vector(15 downto 0) := x"2F";
constant D220: std_logic_vector(15 downto 0) := x"2E";
constant D221: std_logic_vector(15 downto 0) := x"2C";
constant D222: std_logic_vector(15 downto 0) := x"2A";
constant D223: std_logic_vector(15 downto 0) := x"29";
constant D224: std_logic_vector(15 downto 0) := x"27";
constant D225: std_logic_vector(15 downto 0) := x"25";
constant D226: std_logic_vector(15 downto 0) := x"24";
constant D227: std_logic_vector(15 downto 0) := x"22";
constant D228: std_logic_vector(15 downto 0) := x"21";
constant D229: std_logic_vector(15 downto 0) := x"1F";
constant D230: std_logic_vector(15 downto 0) := x"1E";
constant D231: std_logic_vector(15 downto 0) := x"1D";
constant D232: std_logic_vector(15 downto 0) := x"1B";
constant D233: std_logic_vector(15 downto 0) := x"1A";
constant D234: std_logic_vector(15 downto 0) := x"18";
constant D235: std_logic_vector(15 downto 0) := x"17";
constant D236: std_logic_vector(15 downto 0) := x"16";
constant D237: std_logic_vector(15 downto 0) := x"15";
constant D238: std_logic_vector(15 downto 0) := x"13";
constant D239: std_logic_vector(15 downto 0) := x"12";
constant D240: std_logic_vector(15 downto 0) := x"11";
constant D241: std_logic_vector(15 downto 0) := x"10";
constant D242: std_logic_vector(15 downto 0) := x"0F";
constant D243: std_logic_vector(15 downto 0) := x"0E";
constant D244: std_logic_vector(15 downto 0) := x"0D";
constant D245: std_logic_vector(15 downto 0) := x"0C";
constant D246: std_logic_vector(15 downto 0) := x"0B";
constant D247: std_logic_vector(15 downto 0) := x"0A";
constant D248: std_logic_vector(15 downto 0) := x"09";
constant D249: std_logic_vector(15 downto 0) := x"09";
constant D250: std_logic_vector(15 downto 0) := x"08";
constant D251: std_logic_vector(15 downto 0) := x"07";
constant D252: std_logic_vector(15 downto 0) := x"06";
constant D253: std_logic_vector(15 downto 0) := x"06";
constant D254: std_logic_vector(15 downto 0) := x"05";
constant D255: std_logic_vector(15 downto 0) := x"04";
constant D256: std_logic_vector(15 downto 0) := x"04";
constant D257: std_logic_vector(15 downto 0) := x"03";
constant D258: std_logic_vector(15 downto 0) := x"03";
constant D259: std_logic_vector(15 downto 0) := x"02";
constant D260: std_logic_vector(15 downto 0) := x"02";
constant D261: std_logic_vector(15 downto 0) := x"02";
constant D262: std_logic_vector(15 downto 0) := x"01";
constant D263: std_logic_vector(15 downto 0) := x"01";
constant D264: std_logic_vector(15 downto 0) := x"01";
constant D265: std_logic_vector(15 downto 0) := x"00";
constant D266: std_logic_vector(15 downto 0) := x"00";
constant D267: std_logic_vector(15 downto 0) := x"00";
constant D268: std_logic_vector(15 downto 0) := x"00";
constant D269: std_logic_vector(15 downto 0) := x"00";
constant D270: std_logic_vector(15 downto 0) := x"00";
constant D271: std_logic_vector(15 downto 0) := x"00";
constant D272: std_logic_vector(15 downto 0) := x"00";
constant D273: std_logic_vector(15 downto 0) := x"00";
constant D274: std_logic_vector(15 downto 0) := x"00";
constant D275: std_logic_vector(15 downto 0) := x"00";
constant D276: std_logic_vector(15 downto 0) := x"01";
constant D277: std_logic_vector(15 downto 0) := x"01";
constant D278: std_logic_vector(15 downto 0) := x"01";
constant D279: std_logic_vector(15 downto 0) := x"02";
constant D280: std_logic_vector(15 downto 0) := x"02";
constant D281: std_logic_vector(15 downto 0) := x"02";
constant D282: std_logic_vector(15 downto 0) := x"03";
constant D283: std_logic_vector(15 downto 0) := x"03";
constant D284: std_logic_vector(15 downto 0) := x"04";
constant D285: std_logic_vector(15 downto 0) := x"04";
constant D286: std_logic_vector(15 downto 0) := x"05";
constant D287: std_logic_vector(15 downto 0) := x"06";
constant D288: std_logic_vector(15 downto 0) := x"06";
constant D289: std_logic_vector(15 downto 0) := x"07";
constant D290: std_logic_vector(15 downto 0) := x"08";
constant D291: std_logic_vector(15 downto 0) := x"09";
constant D292: std_logic_vector(15 downto 0) := x"09";
constant D293: std_logic_vector(15 downto 0) := x"0A";
constant D294: std_logic_vector(15 downto 0) := x"0B";
constant D295: std_logic_vector(15 downto 0) := x"0C";
constant D296: std_logic_vector(15 downto 0) := x"0D";
constant D297: std_logic_vector(15 downto 0) := x"0E";
constant D298: std_logic_vector(15 downto 0) := x"0F";
constant D299: std_logic_vector(15 downto 0) := x"10";
constant D300: std_logic_vector(15 downto 0) := x"11";
constant D301: std_logic_vector(15 downto 0) := x"12";
constant D302: std_logic_vector(15 downto 0) := x"13";
constant D303: std_logic_vector(15 downto 0) := x"15";
constant D304: std_logic_vector(15 downto 0) := x"16";
constant D305: std_logic_vector(15 downto 0) := x"17";
constant D306: std_logic_vector(15 downto 0) := x"18";
constant D307: std_logic_vector(15 downto 0) := x"1A";
constant D308: std_logic_vector(15 downto 0) := x"1B";
constant D309: std_logic_vector(15 downto 0) := x"1D";
constant D310: std_logic_vector(15 downto 0) := x"1E";
constant D311: std_logic_vector(15 downto 0) := x"1F";
constant D312: std_logic_vector(15 downto 0) := x"21";
constant D313: std_logic_vector(15 downto 0) := x"22";
constant D314: std_logic_vector(15 downto 0) := x"24";
constant D315: std_logic_vector(15 downto 0) := x"25";
constant D316: std_logic_vector(15 downto 0) := x"27";
constant D317: std_logic_vector(15 downto 0) := x"29";
constant D318: std_logic_vector(15 downto 0) := x"2A";
constant D319: std_logic_vector(15 downto 0) := x"2C";
constant D320: std_logic_vector(15 downto 0) := x"2E";
constant D321: std_logic_vector(15 downto 0) := x"2F";
constant D322: std_logic_vector(15 downto 0) := x"31";
constant D323: std_logic_vector(15 downto 0) := x"33";
constant D324: std_logic_vector(15 downto 0) := x"35";
constant D325: std_logic_vector(15 downto 0) := x"37";
constant D326: std_logic_vector(15 downto 0) := x"38";
constant D327: std_logic_vector(15 downto 0) := x"3A";
constant D328: std_logic_vector(15 downto 0) := x"3C";
constant D329: std_logic_vector(15 downto 0) := x"3E";
constant D330: std_logic_vector(15 downto 0) := x"40";
constant D331: std_logic_vector(15 downto 0) := x"42";
constant D332: std_logic_vector(15 downto 0) := x"44";
constant D333: std_logic_vector(15 downto 0) := x"46";
constant D334: std_logic_vector(15 downto 0) := x"48";
constant D335: std_logic_vector(15 downto 0) := x"4A";
constant D336: std_logic_vector(15 downto 0) := x"4C";
constant D337: std_logic_vector(15 downto 0) := x"4E";
constant D338: std_logic_vector(15 downto 0) := x"50";
constant D339: std_logic_vector(15 downto 0) := x"52";
constant D340: std_logic_vector(15 downto 0) := x"54";
constant D341: std_logic_vector(15 downto 0) := x"56";
constant D342: std_logic_vector(15 downto 0) := x"58";
constant D343: std_logic_vector(15 downto 0) := x"5B";
constant D344: std_logic_vector(15 downto 0) := x"5D";
constant D345: std_logic_vector(15 downto 0) := x"5F";
constant D346: std_logic_vector(15 downto 0) := x"61";
constant D347: std_logic_vector(15 downto 0) := x"63";
constant D348: std_logic_vector(15 downto 0) := x"65";
constant D349: std_logic_vector(15 downto 0) := x"68";
constant D350: std_logic_vector(15 downto 0) := x"6A";
constant D351: std_logic_vector(15 downto 0) := x"6C";
constant D352: std_logic_vector(15 downto 0) := x"6E";
constant D353: std_logic_vector(15 downto 0) := x"70";
constant D354: std_logic_vector(15 downto 0) := x"73";
constant D355: std_logic_vector(15 downto 0) := x"75";
constant D356: std_logic_vector(15 downto 0) := x"77";
constant D357: std_logic_vector(15 downto 0) := x"79";
constant D358: std_logic_vector(15 downto 0) := x"7C";
constant D359: std_logic_vector(15 downto 0) := x"7E";
constant D360: std_logic_vector(15 downto 0) := x"80";
type rom_array is array (NATURAL range <>) of STD_LOGIC_VECTOR(15 downto 0);
constant rom: rom_array := (D0,D1,D2,D3,D4,D5,D6,D7,D8,D9,D10,D11,D12,D13,D14,D15,D16,D17,D18,D19,D20,D21,D22,D23,D24,D25,D26,D27,D28,D29,D30,D31,D32,
D33,D34,D35,D36,D37,D38,D39,D40,D41,D42,D43,D44,D45,D46,D47,D48,D49,D50,D51,D52,D53,D54,D55,D56,D57,D58,D59,D60,D61,D62,D63,D64,
D65,D66,D67,D68,D69,D70,D71,D72,D73,D74,D75,D76,D77,D78,D79,D80,D81,D82,D83,D84,D85,D86,D87,D88,D89,D90,D91,D92,D93,D94,D95,D96,
D97,D98,D99,D100,D101,D102,D103,D104,D105,D106,D107,D108,D109,D110,D111,D112,D113,D114,D115,D116,D117,D118,D119,D120,D121,D122,D123,D124,D125,D126,D127,D128,
D129,D130,D131,D132,D133,D134,D135,D136,D137,D138,D139,D140,D141,D142,D143,D144,D145,D146,D147,D148,D149,D150,D151,D152,D153,D154,D155,D156,D157,D158,D159,D160,
D161,D162,D163,D164,D165,D166,D167,D168,D169,D170,D171,D172,D173,D174,D175,D176,D177,D178,D179,D180,D181,D182,D183,D184,D185,D186,D187,D188,D189,D190,D191,D192,
D193,D194,D195,D196,D197,D198,D199,D200,D201,D202,D203,D204,D205,D206,D207,D208,D209,D210,D211,D212,D213,D214,D215,D216,D217,D218,D219,D220,D221,D222,D223,D224,
D225,D226,D227,D228,D229,D230,D231,D232,D233,D234,D235,D236,D237,D238,D239,D240,D241,D242,D243,D244,D245,D246,D247,D248,D249,D250,D251,D252,D253,D254,D255,D256,
D257,D258,D259,D260,D261,D262,D263,D264,D265,D266,D267,D268,D269,D270,D271,D272,D273,D274,D275,D276,D277,D278,D279,D280,D281,D282,D283,D284,D285,D286,D287,D288,
D289,D290,D291,D292,D293,D294,D295,D296,D297,D298,D299,D300,D301,D302,D303,D304,D305,D306,D307,D308,D309,D310,D311,D312,D313,D314,D315,D316,D317,D318,D319,D320,
D321,D322,D323,D324,D325,D326,D327,D328,D329,D330,D331,D332,D333,D334,D335,D336,D337,D338,D339,D340,D341,D342,D343,D344,D345,D346,D347,D348,D349,D350,D351,D352,
D353,D354,D355,D356,D357,D358,D359,D360,);
begin
process(clk)
variable j: integer;
begin
if(rising_edge(clk)) then  j := conv_integer(dir);
dataout <= rom(j); 
j<= j+1
if(j=180) then
j<=0;
end if;
end if;
end process;
end Behavioral;

