library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
entity TriangleWave is
port (clksen :in  std_logic;
dataout : out std_logic_vector(15 downto 0);
);
end TriangleWave;
architecture Behavioral of TriangleWave is


constant dato0: std_logic_vector(15 downto 0) := x"80";
constant dato1: std_logic_vector(15 downto 0) := x"81";
constant dato2: std_logic_vector(15 downto 0) := x"83";
constant dato3: std_logic_vector(15 downto 0) := x"84";
constant dato4: std_logic_vector(15 downto 0) := x"86";
constant dato5: std_logic_vector(15 downto 0) := x"87";
constant dato6: std_logic_vector(15 downto 0) := x"88";
constant dato7: std_logic_vector(15 downto 0) := x"8A";
constant dato8: std_logic_vector(15 downto 0) := x"8B";
constant dato9: std_logic_vector(15 downto 0) := x"8D";
constant dato10: std_logic_vector(15 downto 0) := x"8E";
constant dato11: std_logic_vector(15 downto 0) := x"90";
constant dato12: std_logic_vector(15 downto 0) := x"91";
constant dato13: std_logic_vector(15 downto 0) := x"92";
constant dato14: std_logic_vector(15 downto 0) := x"94";
constant dato15: std_logic_vector(15 downto 0) := x"95";
constant dato16: std_logic_vector(15 downto 0) := x"97";
constant dato17: std_logic_vector(15 downto 0) := x"98";
constant dato18: std_logic_vector(15 downto 0) := x"99";
constant dato19: std_logic_vector(15 downto 0) := x"9B";
constant dato20: std_logic_vector(15 downto 0) := x"9C";
constant dato21: std_logic_vector(15 downto 0) := x"9E";
constant dato22: std_logic_vector(15 downto 0) := x"9F";
constant dato23: std_logic_vector(15 downto 0) := x"A0";
constant dato24: std_logic_vector(15 downto 0) := x"A2";
constant dato25: std_logic_vector(15 downto 0) := x"A3";
constant dato26: std_logic_vector(15 downto 0) := x"A5";
constant dato27: std_logic_vector(15 downto 0) := x"A6";
constant dato28: std_logic_vector(15 downto 0) := x"A7";
constant dato29: std_logic_vector(15 downto 0) := x"A9";
constant dato30: std_logic_vector(15 downto 0) := x"AA";
constant dato31: std_logic_vector(15 downto 0) := x"AC";
constant dato32: std_logic_vector(15 downto 0) := x"AD";
constant dato33: std_logic_vector(15 downto 0) := x"AF";
constant dato34: std_logic_vector(15 downto 0) := x"B0";
constant dato35: std_logic_vector(15 downto 0) := x"B1";
constant dato36: std_logic_vector(15 downto 0) := x"B3";
constant dato37: std_logic_vector(15 downto 0) := x"B4";
constant dato38: std_logic_vector(15 downto 0) := x"B6";
constant dato39: std_logic_vector(15 downto 0) := x"B7";
constant dato40: std_logic_vector(15 downto 0) := x"B8";
constant dato41: std_logic_vector(15 downto 0) := x"BA";
constant dato42: std_logic_vector(15 downto 0) := x"BB";
constant dato43: std_logic_vector(15 downto 0) := x"BD";
constant dato44: std_logic_vector(15 downto 0) := x"BE";
constant dato45: std_logic_vector(15 downto 0) := x"BF";
constant dato46: std_logic_vector(15 downto 0) := x"C1";
constant dato47: std_logic_vector(15 downto 0) := x"C2";
constant dato48: std_logic_vector(15 downto 0) := x"C4";
constant dato49: std_logic_vector(15 downto 0) := x"C5";
constant dato50: std_logic_vector(15 downto 0) := x"C7";
constant dato51: std_logic_vector(15 downto 0) := x"C8";
constant dato52: std_logic_vector(15 downto 0) := x"C9";
constant dato53: std_logic_vector(15 downto 0) := x"CB";
constant dato54: std_logic_vector(15 downto 0) := x"CC";
constant dato55: std_logic_vector(15 downto 0) := x"CE";
constant dato56: std_logic_vector(15 downto 0) := x"CF";
constant dato57: std_logic_vector(15 downto 0) := x"D0";
constant dato58: std_logic_vector(15 downto 0) := x"D2";
constant dato59: std_logic_vector(15 downto 0) := x"D3";
constant dato60: std_logic_vector(15 downto 0) := x"D5";
constant dato61: std_logic_vector(15 downto 0) := x"D6";
constant dato62: std_logic_vector(15 downto 0) := x"D7";
constant dato63: std_logic_vector(15 downto 0) := x"D9";
constant dato64: std_logic_vector(15 downto 0) := x"DA";
constant dato65: std_logic_vector(15 downto 0) := x"DC";
constant dato66: std_logic_vector(15 downto 0) := x"DD";
constant dato67: std_logic_vector(15 downto 0) := x"DE";
constant dato68: std_logic_vector(15 downto 0) := x"E0";
constant dato69: std_logic_vector(15 downto 0) := x"E1";
constant dato70: std_logic_vector(15 downto 0) := x"E3";
constant dato71: std_logic_vector(15 downto 0) := x"E4";
constant dato72: std_logic_vector(15 downto 0) := x"E6";
constant dato73: std_logic_vector(15 downto 0) := x"E7";
constant dato74: std_logic_vector(15 downto 0) := x"E8";
constant dato75: std_logic_vector(15 downto 0) := x"EA";
constant dato76: std_logic_vector(15 downto 0) := x"EB";
constant dato77: std_logic_vector(15 downto 0) := x"ED";
constant dato78: std_logic_vector(15 downto 0) := x"EE";
constant dato79: std_logic_vector(15 downto 0) := x"EF";
constant dato80: std_logic_vector(15 downto 0) := x"F1";
constant dato81: std_logic_vector(15 downto 0) := x"F2";
constant dato82: std_logic_vector(15 downto 0) := x"F4";
constant dato83: std_logic_vector(15 downto 0) := x"F5";
constant dato84: std_logic_vector(15 downto 0) := x"F6";
constant dato85: std_logic_vector(15 downto 0) := x"F8";
constant dato86: std_logic_vector(15 downto 0) := x"F9";
constant dato87: std_logic_vector(15 downto 0) := x"FB";
constant dato88: std_logic_vector(15 downto 0) := x"FC";
constant dato89: std_logic_vector(15 downto 0) := x"FD";
constant dato90: std_logic_vector(15 downto 0) := x"FF";
constant dato91: std_logic_vector(15 downto 0) := x"FF";
constant dato92: std_logic_vector(15 downto 0) := x"FD";
constant dato93: std_logic_vector(15 downto 0) := x"FC";
constant dato94: std_logic_vector(15 downto 0) := x"FA";
constant dato95: std_logic_vector(15 downto 0) := x"F9";
constant dato96: std_logic_vector(15 downto 0) := x"F8";
constant dato97: std_logic_vector(15 downto 0) := x"F6";
constant dato98: std_logic_vector(15 downto 0) := x"F5";
constant dato99: std_logic_vector(15 downto 0) := x"F3";
constant dato100: std_logic_vector(15 downto 0) := x"F2";
constant dato101: std_logic_vector(15 downto 0) := x"F1";
constant dato102: std_logic_vector(15 downto 0) := x"EF";
constant dato103: std_logic_vector(15 downto 0) := x"EE";
constant dato104: std_logic_vector(15 downto 0) := x"EC";
constant dato105: std_logic_vector(15 downto 0) := x"EB";
constant dato106: std_logic_vector(15 downto 0) := x"EA";
constant dato107: std_logic_vector(15 downto 0) := x"E8";
constant dato108: std_logic_vector(15 downto 0) := x"E7";
constant dato109: std_logic_vector(15 downto 0) := x"E5";
constant dato110: std_logic_vector(15 downto 0) := x"E4";
constant dato111: std_logic_vector(15 downto 0) := x"E2";
constant dato112: std_logic_vector(15 downto 0) := x"E1";
constant dato113: std_logic_vector(15 downto 0) := x"E0";
constant dato114: std_logic_vector(15 downto 0) := x"DE";
constant dato115: std_logic_vector(15 downto 0) := x"DD";
constant dato116: std_logic_vector(15 downto 0) := x"DB";
constant dato117: std_logic_vector(15 downto 0) := x"DA";
constant dato118: std_logic_vector(15 downto 0) := x"D9";
constant dato119: std_logic_vector(15 downto 0) := x"D7";
constant dato120: std_logic_vector(15 downto 0) := x"D6";
constant dato121: std_logic_vector(15 downto 0) := x"D4";
constant dato122: std_logic_vector(15 downto 0) := x"D3";
constant dato123: std_logic_vector(15 downto 0) := x"D2";
constant dato124: std_logic_vector(15 downto 0) := x"D0";
constant dato125: std_logic_vector(15 downto 0) := x"CF";
constant dato126: std_logic_vector(15 downto 0) := x"CD";
constant dato127: std_logic_vector(15 downto 0) := x"CC";
constant dato128: std_logic_vector(15 downto 0) := x"CB";
constant dato129: std_logic_vector(15 downto 0) := x"C9";
constant dato130: std_logic_vector(15 downto 0) := x"C8";
constant dato131: std_logic_vector(15 downto 0) := x"C6";
constant dato132: std_logic_vector(15 downto 0) := x"C5";
constant dato133: std_logic_vector(15 downto 0) := x"C3";
constant dato134: std_logic_vector(15 downto 0) := x"C2";
constant dato135: std_logic_vector(15 downto 0) := x"C1";
constant dato136: std_logic_vector(15 downto 0) := x"BF";
constant dato137: std_logic_vector(15 downto 0) := x"BE";
constant dato138: std_logic_vector(15 downto 0) := x"BC";
constant dato139: std_logic_vector(15 downto 0) := x"BB";
constant dato140: std_logic_vector(15 downto 0) := x"BA";
constant dato141: std_logic_vector(15 downto 0) := x"B8";
constant dato142: std_logic_vector(15 downto 0) := x"B7";
constant dato143: std_logic_vector(15 downto 0) := x"B5";
constant dato144: std_logic_vector(15 downto 0) := x"B4";
constant dato145: std_logic_vector(15 downto 0) := x"B3";
constant dato146: std_logic_vector(15 downto 0) := x"B1";
constant dato147: std_logic_vector(15 downto 0) := x"B0";
constant dato148: std_logic_vector(15 downto 0) := x"AE";
constant dato149: std_logic_vector(15 downto 0) := x"AD";
constant dato150: std_logic_vector(15 downto 0) := x"AB";
constant dato151: std_logic_vector(15 downto 0) := x"AA";
constant dato152: std_logic_vector(15 downto 0) := x"A9";
constant dato153: std_logic_vector(15 downto 0) := x"A7";
constant dato154: std_logic_vector(15 downto 0) := x"A6";
constant dato155: std_logic_vector(15 downto 0) := x"A4";
constant dato156: std_logic_vector(15 downto 0) := x"A3";
constant dato157: std_logic_vector(15 downto 0) := x"A2";
constant dato158: std_logic_vector(15 downto 0) := x"A0";
constant dato159: std_logic_vector(15 downto 0) := x"9F";
constant dato160: std_logic_vector(15 downto 0) := x"9D";
constant dato161: std_logic_vector(15 downto 0) := x"9C";
constant dato162: std_logic_vector(15 downto 0) := x"9B";
constant dato163: std_logic_vector(15 downto 0) := x"99";
constant dato164: std_logic_vector(15 downto 0) := x"98";
constant dato165: std_logic_vector(15 downto 0) := x"96";
constant dato166: std_logic_vector(15 downto 0) := x"95";
constant dato167: std_logic_vector(15 downto 0) := x"94";
constant dato168: std_logic_vector(15 downto 0) := x"92";
constant dato169: std_logic_vector(15 downto 0) := x"91";
constant dato170: std_logic_vector(15 downto 0) := x"8F";
constant dato171: std_logic_vector(15 downto 0) := x"8E";
constant dato172: std_logic_vector(15 downto 0) := x"8C";
constant dato173: std_logic_vector(15 downto 0) := x"8B";
constant dato174: std_logic_vector(15 downto 0) := x"8A";
constant dato175: std_logic_vector(15 downto 0) := x"88";
constant dato176: std_logic_vector(15 downto 0) := x"87";
constant dato177: std_logic_vector(15 downto 0) := x"85";
constant dato178: std_logic_vector(15 downto 0) := x"84";
constant dato179: std_logic_vector(15 downto 0) := x"83";
constant dato180: std_logic_vector(15 downto 0) := x"81";
constant dato181: std_logic_vector(15 downto 0) := x"80";
constant dato182: std_logic_vector(15 downto 0) := x"7E";
constant dato183: std_logic_vector(15 downto 0) := x"7D";
constant dato184: std_logic_vector(15 downto 0) := x"7C";
constant dato185: std_logic_vector(15 downto 0) := x"7A";
constant dato186: std_logic_vector(15 downto 0) := x"79";
constant dato187: std_logic_vector(15 downto 0) := x"77";
constant dato188: std_logic_vector(15 downto 0) := x"76";
constant dato189: std_logic_vector(15 downto 0) := x"75";
constant dato190: std_logic_vector(15 downto 0) := x"73";
constant dato191: std_logic_vector(15 downto 0) := x"72";
constant dato192: std_logic_vector(15 downto 0) := x"70";
constant dato193: std_logic_vector(15 downto 0) := x"6F";
constant dato194: std_logic_vector(15 downto 0) := x"6D";
constant dato195: std_logic_vector(15 downto 0) := x"6C";
constant dato196: std_logic_vector(15 downto 0) := x"6B";
constant dato197: std_logic_vector(15 downto 0) := x"69";
constant dato198: std_logic_vector(15 downto 0) := x"68";
constant dato199: std_logic_vector(15 downto 0) := x"66";
constant dato200: std_logic_vector(15 downto 0) := x"65";
constant dato201: std_logic_vector(15 downto 0) := x"64";
constant dato202: std_logic_vector(15 downto 0) := x"62";
constant dato203: std_logic_vector(15 downto 0) := x"61";
constant dato204: std_logic_vector(15 downto 0) := x"5F";
constant dato205: std_logic_vector(15 downto 0) := x"5E";
constant dato206: std_logic_vector(15 downto 0) := x"5D";
constant dato207: std_logic_vector(15 downto 0) := x"5B";
constant dato208: std_logic_vector(15 downto 0) := x"5A";
constant dato209: std_logic_vector(15 downto 0) := x"58";
constant dato210: std_logic_vector(15 downto 0) := x"57";
constant dato211: std_logic_vector(15 downto 0) := x"55";
constant dato212: std_logic_vector(15 downto 0) := x"54";
constant dato213: std_logic_vector(15 downto 0) := x"53";
constant dato214: std_logic_vector(15 downto 0) := x"51";
constant dato215: std_logic_vector(15 downto 0) := x"50";
constant dato216: std_logic_vector(15 downto 0) := x"4E";
constant dato217: std_logic_vector(15 downto 0) := x"4D";
constant dato218: std_logic_vector(15 downto 0) := x"4C";
constant dato219: std_logic_vector(15 downto 0) := x"4A";
constant dato220: std_logic_vector(15 downto 0) := x"49";
constant dato221: std_logic_vector(15 downto 0) := x"47";
constant dato222: std_logic_vector(15 downto 0) := x"46";
constant dato223: std_logic_vector(15 downto 0) := x"45";
constant dato224: std_logic_vector(15 downto 0) := x"43";
constant dato225: std_logic_vector(15 downto 0) := x"42";
constant dato226: std_logic_vector(15 downto 0) := x"40";
constant dato227: std_logic_vector(15 downto 0) := x"3F";
constant dato228: std_logic_vector(15 downto 0) := x"3E";
constant dato229: std_logic_vector(15 downto 0) := x"3C";
constant dato230: std_logic_vector(15 downto 0) := x"3B";
constant dato231: std_logic_vector(15 downto 0) := x"39";
constant dato232: std_logic_vector(15 downto 0) := x"38";
constant dato233: std_logic_vector(15 downto 0) := x"36";
constant dato234: std_logic_vector(15 downto 0) := x"35";
constant dato235: std_logic_vector(15 downto 0) := x"34";
constant dato236: std_logic_vector(15 downto 0) := x"32";
constant dato237: std_logic_vector(15 downto 0) := x"31";
constant dato238: std_logic_vector(15 downto 0) := x"2F";
constant dato239: std_logic_vector(15 downto 0) := x"2E";
constant dato240: std_logic_vector(15 downto 0) := x"2D";
constant dato241: std_logic_vector(15 downto 0) := x"2B";
constant dato242: std_logic_vector(15 downto 0) := x"2A";
constant dato243: std_logic_vector(15 downto 0) := x"28";
constant dato244: std_logic_vector(15 downto 0) := x"27";
constant dato245: std_logic_vector(15 downto 0) := x"26";
constant dato246: std_logic_vector(15 downto 0) := x"24";
constant dato247: std_logic_vector(15 downto 0) := x"23";
constant dato248: std_logic_vector(15 downto 0) := x"21";
constant dato249: std_logic_vector(15 downto 0) := x"20";
constant dato250: std_logic_vector(15 downto 0) := x"1E";
constant dato251: std_logic_vector(15 downto 0) := x"1D";
constant dato252: std_logic_vector(15 downto 0) := x"1C";
constant dato253: std_logic_vector(15 downto 0) := x"1A";
constant dato254: std_logic_vector(15 downto 0) := x"19";
constant dato255: std_logic_vector(15 downto 0) := x"17";
constant dato256: std_logic_vector(15 downto 0) := x"16";
constant dato257: std_logic_vector(15 downto 0) := x"15";
constant dato258: std_logic_vector(15 downto 0) := x"13";
constant dato259: std_logic_vector(15 downto 0) := x"12";
constant dato260: std_logic_vector(15 downto 0) := x"10";
constant dato261: std_logic_vector(15 downto 0) := x"0F";
constant dato262: std_logic_vector(15 downto 0) := x"0E";
constant dato263: std_logic_vector(15 downto 0) := x"0C";
constant dato264: std_logic_vector(15 downto 0) := x"0B";
constant dato265: std_logic_vector(15 downto 0) := x"09";
constant dato266: std_logic_vector(15 downto 0) := x"08";
constant dato267: std_logic_vector(15 downto 0) := x"07";
constant dato268: std_logic_vector(15 downto 0) := x"05";
constant dato269: std_logic_vector(15 downto 0) := x"04";
constant dato270: std_logic_vector(15 downto 0) := x"02";
constant dato271: std_logic_vector(15 downto 0) := x"02";
constant dato272: std_logic_vector(15 downto 0) := x"04";
constant dato273: std_logic_vector(15 downto 0) := x"05";
constant dato274: std_logic_vector(15 downto 0) := x"06";
constant dato275: std_logic_vector(15 downto 0) := x"08";
constant dato276: std_logic_vector(15 downto 0) := x"09";
constant dato277: std_logic_vector(15 downto 0) := x"0B";
constant dato278: std_logic_vector(15 downto 0) := x"0C";
constant dato279: std_logic_vector(15 downto 0) := x"0D";
constant dato280: std_logic_vector(15 downto 0) := x"0F";
constant dato281: std_logic_vector(15 downto 0) := x"10";
constant dato282: std_logic_vector(15 downto 0) := x"12";
constant dato283: std_logic_vector(15 downto 0) := x"13";
constant dato284: std_logic_vector(15 downto 0) := x"14";
constant dato285: std_logic_vector(15 downto 0) := x"16";
constant dato286: std_logic_vector(15 downto 0) := x"17";
constant dato287: std_logic_vector(15 downto 0) := x"19";
constant dato288: std_logic_vector(15 downto 0) := x"1A";
constant dato289: std_logic_vector(15 downto 0) := x"1B";
constant dato290: std_logic_vector(15 downto 0) := x"1D";
constant dato291: std_logic_vector(15 downto 0) := x"1E";
constant dato292: std_logic_vector(15 downto 0) := x"20";
constant dato293: std_logic_vector(15 downto 0) := x"21";
constant dato294: std_logic_vector(15 downto 0) := x"23";
constant dato295: std_logic_vector(15 downto 0) := x"24";
constant dato296: std_logic_vector(15 downto 0) := x"25";
constant dato297: std_logic_vector(15 downto 0) := x"27";
constant dato298: std_logic_vector(15 downto 0) := x"28";
constant dato299: std_logic_vector(15 downto 0) := x"2A";
constant dato300: std_logic_vector(15 downto 0) := x"2B";
constant dato301: std_logic_vector(15 downto 0) := x"2C";
constant dato302: std_logic_vector(15 downto 0) := x"2E";
constant dato303: std_logic_vector(15 downto 0) := x"2F";
constant dato304: std_logic_vector(15 downto 0) := x"31";
constant dato305: std_logic_vector(15 downto 0) := x"32";
constant dato306: std_logic_vector(15 downto 0) := x"33";
constant dato307: std_logic_vector(15 downto 0) := x"35";
constant dato308: std_logic_vector(15 downto 0) := x"36";
constant dato309: std_logic_vector(15 downto 0) := x"38";
constant dato310: std_logic_vector(15 downto 0) := x"39";
constant dato311: std_logic_vector(15 downto 0) := x"3B";
constant dato312: std_logic_vector(15 downto 0) := x"3C";
constant dato313: std_logic_vector(15 downto 0) := x"3D";
constant dato314: std_logic_vector(15 downto 0) := x"3F";
constant dato315: std_logic_vector(15 downto 0) := x"40";
constant dato316: std_logic_vector(15 downto 0) := x"42";
constant dato317: std_logic_vector(15 downto 0) := x"43";
constant dato318: std_logic_vector(15 downto 0) := x"44";
constant dato319: std_logic_vector(15 downto 0) := x"46";
constant dato320: std_logic_vector(15 downto 0) := x"47";
constant dato321: std_logic_vector(15 downto 0) := x"49";
constant dato322: std_logic_vector(15 downto 0) := x"4A";
constant dato323: std_logic_vector(15 downto 0) := x"4B";
constant dato324: std_logic_vector(15 downto 0) := x"4D";
constant dato325: std_logic_vector(15 downto 0) := x"4E";
constant dato326: std_logic_vector(15 downto 0) := x"50";
constant dato327: std_logic_vector(15 downto 0) := x"51";
constant dato328: std_logic_vector(15 downto 0) := x"52";
constant dato329: std_logic_vector(15 downto 0) := x"54";
constant dato330: std_logic_vector(15 downto 0) := x"55";
constant dato331: std_logic_vector(15 downto 0) := x"57";
constant dato332: std_logic_vector(15 downto 0) := x"58";
constant dato333: std_logic_vector(15 downto 0) := x"5A";
constant dato334: std_logic_vector(15 downto 0) := x"5B";
constant dato335: std_logic_vector(15 downto 0) := x"5C";
constant dato336: std_logic_vector(15 downto 0) := x"5E";
constant dato337: std_logic_vector(15 downto 0) := x"5F";
constant dato338: std_logic_vector(15 downto 0) := x"61";
constant dato339: std_logic_vector(15 downto 0) := x"62";
constant dato340: std_logic_vector(15 downto 0) := x"63";
constant dato341: std_logic_vector(15 downto 0) := x"65";
constant dato342: std_logic_vector(15 downto 0) := x"66";
constant dato343: std_logic_vector(15 downto 0) := x"68";
constant dato344: std_logic_vector(15 downto 0) := x"69";
constant dato345: std_logic_vector(15 downto 0) := x"6A";
constant dato346: std_logic_vector(15 downto 0) := x"6C";
constant dato347: std_logic_vector(15 downto 0) := x"6D";
constant dato348: std_logic_vector(15 downto 0) := x"6F";
constant dato349: std_logic_vector(15 downto 0) := x"70";
constant dato350: std_logic_vector(15 downto 0) := x"72";
constant dato351: std_logic_vector(15 downto 0) := x"73";
constant dato352: std_logic_vector(15 downto 0) := x"74";
constant dato353: std_logic_vector(15 downto 0) := x"76";
constant dato354: std_logic_vector(15 downto 0) := x"77";
constant dato355: std_logic_vector(15 downto 0) := x"79";
constant dato356: std_logic_vector(15 downto 0) := x"7A";
constant dato357: std_logic_vector(15 downto 0) := x"7B";
constant dato358: std_logic_vector(15 downto 0) := x"7D";
constant dato359: std_logic_vector(15 downto 0) := x"7E";
constant dato360: std_logic_vector(15 downto 0) := x"80";
type rom_array is array (NATURAL range <>) of STD_LOGIC_VECTOR(15 downto 0);
constant rom: rom_array := (D0,D1,D2,D3,D4,D5,D6,D7,D8,D9,D10,D11,D12,D13,D14,D15,D16,D17,D18,D19,D20,D21,D22,D23,D24,D25,D26,D27,D28,D29,D30,D31,D32,
D33,D34,D35,D36,D37,D38,D39,D40,D41,D42,D43,D44,D45,D46,D47,D48,D49,D50,D51,D52,D53,D54,D55,D56,D57,D58,D59,D60,D61,D62,D63,D64,
D65,D66,D67,D68,D69,D70,D71,D72,D73,D74,D75,D76,D77,D78,D79,D80,D81,D82,D83,D84,D85,D86,D87,D88,D89,D90,D91,D92,D93,D94,D95,D96,
D97,D98,D99,D100,D101,D102,D103,D104,D105,D106,D107,D108,D109,D110,D111,D112,D113,D114,D115,D116,D117,D118,D119,D120,D121,D122,D123,D124,D125,D126,D127,D128,
D129,D130,D131,D132,D133,D134,D135,D136,D137,D138,D139,D140,D141,D142,D143,D144,D145,D146,D147,D148,D149,D150,D151,D152,D153,D154,D155,D156,D157,D158,D159,D160,
D161,D162,D163,D164,D165,D166,D167,D168,D169,D170,D171,D172,D173,D174,D175,D176,D177,D178,D179,D180,D181,D182,D183,D184,D185,D186,D187,D188,D189,D190,D191,D192,
D193,D194,D195,D196,D197,D198,D199,D200,D201,D202,D203,D204,D205,D206,D207,D208,D209,D210,D211,D212,D213,D214,D215,D216,D217,D218,D219,D220,D221,D222,D223,D224,
D225,D226,D227,D228,D229,D230,D231,D232,D233,D234,D235,D236,D237,D238,D239,D240,D241,D242,D243,D244,D245,D246,D247,D248,D249,D250,D251,D252,D253,D254,D255,D256,
D257,D258,D259,D260,D261,D262,D263,D264,D265,D266,D267,D268,D269,D270,D271,D272,D273,D274,D275,D276,D277,D278,D279,D280,D281,D282,D283,D284,D285,D286,D287,D288,
D289,D290,D291,D292,D293,D294,D295,D296,D297,D298,D299,D300,D301,D302,D303,D304,D305,D306,D307,D308,D309,D310,D311,D312,D313,D314,D315,D316,D317,D318,D319,D320,
D321,D322,D323,D324,D325,D326,D327,D328,D329,D330,D331,D332,D333,D334,D335,D336,D337,D338,D339,D340,D341,D342,D343,D344,D345,D346,D347,D348,D349,D350,D351,D352,
D353,D354,D355,D356,D357,D358,D359,D360,);
begin
process(clksen)
variable j: integer;
begin
if(rising_edge(clk)) then  j := conv_integer(dir);
dataout <= rom(j); 
j<= j+1
if(j=180) then
j<=0;
end if;
end if;
end process;
end Behavioral;

