library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DigitalControlledOsc is
end DigitalControlledOsc;

architecture Behavioral of DigitalControlledOsc is

begin


end Behavioral;

