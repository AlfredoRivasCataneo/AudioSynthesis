library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DigitalControlledAmp is
end DigitalControlledAmp;

architecture Behavioral of DigitalControlledAmp is

begin


end Behavioral;

